module F1 (f , j , VV1V); 
input f , j;
output VV1V;
or f0 (VV1V , f , j);
endmodule