module F2 (h , f , VV2V); 
input h , f;
output VV2V;
or f0 (VV2V , h , f);
endmodule