module F4 (k , e , VV4V); 
input k , e;
output VV4V;
xor f0 (VV4V , k , e);
endmodule